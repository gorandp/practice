library IEEE;

entity